<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-4.125,10.125,56.275,-56.075</PageViewport>
<gate>
<ID>2</ID>
<type>GA_LED</type>
<position>19.5,-19</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>GA_LED</type>
<position>19.5,-7.5</position>
<input>
<ID>N_in3</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>12,-7.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>4.5,-9</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>4.5,-6.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_OR2</type>
<position>12.5,-19</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>4.5,-18</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>4.5,-21</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>BA_NAND2</type>
<position>32.5,-7</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>24,-6</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>24,-9.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>39.5,-7.5</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AI_XOR2</type>
<position>11.5,-32.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>4.5,-31</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>4.5,-33.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>19.5,-32.5</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_INVERTER</type>
<position>14.5,-46.5</position>
<input>
<ID>IN_0</ID>15 </input>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>9,-46.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>20.5,-46.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AO_XNOR2</type>
<position>31.5,-32.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>24,-31.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>24,-34.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>37.5,-32.5</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>BE_NOR2</type>
<position>31,-20</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>37.5,-20</position>
<input>
<ID>N_in0</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>23.5,-18.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>23.5,-21</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>11.5,-2.5</position>
<gparam>LABEL_TEXT AND GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>31.5,-2</position>
<gparam>LABEL_TEXT NAND GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>10,-14.5</position>
<gparam>LABEL_TEXT OR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>30.5,-14.5</position>
<gparam>LABEL_TEXT NOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>11,-27.5</position>
<gparam>LABEL_TEXT XOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_LABEL</type>
<position>31.5,-27.5</position>
<gparam>LABEL_TEXT XNOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>13,-41</position>
<gparam>LABEL_TEXT NOT GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-7.5,19.5,-6.5</points>
<connection>
<GID>4</GID>
<name>N_in3</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-7.5,19.5,-7.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6.5,-6.5,9,-6.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-9,7.5,-8.5</points>
<intersection>-9 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,-8.5,9,-8.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-9,7.5,-9</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,-19,18.5,-19</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>2</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-21,8,-20</points>
<intersection>-21 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-20,9.5,-20</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6.5,-21,8,-21</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6.5,-18,9.5,-18</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-6,29.5,-6</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-9.5,27.5,-8</points>
<intersection>-9.5 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-8,29.5,-8</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-9.5,27.5,-9.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-7,38.5,-7</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>38.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>38.5,-7.5,38.5,-7</points>
<connection>
<GID>24</GID>
<name>N_in0</name></connection>
<intersection>-7 1</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6.5,-33.5,8.5,-33.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<connection>
<GID>26</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6.5,-31.5,8.5,-31.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>6.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>6.5,-31.5,6.5,-31</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-32.5,18.5,-32.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>32</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>13</ID>
<points>11,-46.5,11.5,-46.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-46.5,19.5,-46.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<connection>
<GID>38</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-34.5,27,-33.5</points>
<intersection>-34.5 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-33.5,28.5,-33.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-34.5,27,-34.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-31.5,28.5,-31.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-32.5,36.5,-32.5</points>
<connection>
<GID>48</GID>
<name>N_in0</name></connection>
<connection>
<GID>40</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-20,36.5,-20</points>
<connection>
<GID>52</GID>
<name>N_in0</name></connection>
<connection>
<GID>50</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-19,26.5,-18.5</points>
<intersection>-19 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-19,28,-19</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-18.5,26.5,-18.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-21,28,-21</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<connection>
<GID>50</GID>
<name>IN_1</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-51.0504,77.2043,56.3273,-40.4846</PageViewport>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>-31.5,42</position>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>-31.5,34.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_INVERTER</type>
<position>-24,37.5</position>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>66</ID>
<type>AE_OR2</type>
<position>1,41</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_AND2</type>
<position>-15.5,36.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_AND2</type>
<position>-15,29</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>-31.5,28</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AI_XOR2</type>
<position>10.5,34.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>GA_LED</type>
<position>16,34.5</position>
<input>
<ID>N_in0</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>-18.5,44.5</position>
<gparam>LABEL_TEXT 32.</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_AND2</type>
<position>-11,10</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AI_XOR2</type>
<position>-19,5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>-31.5,5</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>90</ID>
<type>AA_TOGGLE</type>
<position>-31.5,-1</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_AND2</type>
<position>-17.5,-7</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_TOGGLE</type>
<position>-32,-8</position>
<output>
<ID>OUT_0</ID>36 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>98</ID>
<type>BA_NAND2</type>
<position>-7.5,-12</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AO_XNOR2</type>
<position>-4.5,-1</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AI_XOR2</type>
<position>5,-7</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AE_OR2</type>
<position>12.5,7</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>GA_LED</type>
<position>18,7</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>-2,14</position>
<gparam>LABEL_TEXT 34.</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29.5,42,-2,42</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-27 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27,37.5,-27,42</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>42 1</intersection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-21,37.5,-18.5,37.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>-20 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-20,30,-20,37.5</points>
<intersection>30 3</intersection>
<intersection>37.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-20,30,-18,30</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-20 2</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24,34.5,-24,35.5</points>
<intersection>34.5 2</intersection>
<intersection>35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,35.5,-18.5,35.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>-24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,34.5,-24,34.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>-24 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-29.5,28,-18,28</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<intersection>-18 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-18,28,-18,28</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>28 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-7.5,36.5,-7.5,40</points>
<intersection>36.5 2</intersection>
<intersection>40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-7.5,40,-2,40</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>-7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12.5,36.5,-7.5,36.5</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>-7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,29,-2.5,33.5</points>
<intersection>29 2</intersection>
<intersection>33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,33.5,7.5,33.5</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>-2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-12,29,-2.5,29</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>-2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>5.5,35.5,5.5,41</points>
<intersection>35.5 1</intersection>
<intersection>41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,35.5,7.5,35.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4,41,5.5,41</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,34.5,15,34.5</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<connection>
<GID>76</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,6,-26.5,11</points>
<intersection>6 1</intersection>
<intersection>11 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,6,-22,6</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>-29.5 6</intersection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-26.5,11,-14,11</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-29.5,5,-29.5,6</points>
<intersection>5 9</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-29.5,5,-29.5,5</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>-29.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-24.5,-6,-24.5,4</points>
<intersection>-6 3</intersection>
<intersection>-1 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24.5,4,-22,4</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>-24.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29.5,-1,-24.5,-1</points>
<connection>
<GID>90</GID>
<name>OUT_0</name></connection>
<intersection>-24.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-24.5,-6,-20.5,-6</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>-24.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30,-8,-20.5,-8</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>-26 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-26,-13,-26,-8</points>
<intersection>-13 4</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-26,-13,-10.5,-13</points>
<connection>
<GID>98</GID>
<name>IN_1</name></connection>
<intersection>-26 3</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-11,-12.5,-2</points>
<intersection>-11 1</intersection>
<intersection>-7 2</intersection>
<intersection>-2 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-12.5,-11,-10.5,-11</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-14.5,-7,-12.5,-7</points>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-12.5,-2,-7.5,-2</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>-12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,0,-14,9</points>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>0 2</intersection>
<intersection>5 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14,0,-7.5,0</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-16,5,-14,5</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,-6,1.5,-1</points>
<intersection>-6 3</intersection>
<intersection>-1 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,-1,1.5,-1</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<intersection>1.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>1.5,-6,2,-6</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-12,0.5,-8</points>
<intersection>-12 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-8,2,-8</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4.5,-12,0.5,-12</points>
<connection>
<GID>98</GID>
<name>OUT</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-7,7.5,6</points>
<intersection>-7 2</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7.5,6,9.5,6</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>7.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-7,8,-7</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1,8,1,10</points>
<intersection>8 1</intersection>
<intersection>10 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,8,9.5,8</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>1 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,10,1,10</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<intersection>1 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15.5,7,17,7</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<connection>
<GID>110</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,0,60.4,-66.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,60.4,-66.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,60.4,-66.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,60.4,-66.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,60.4,-66.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,60.4,-66.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,60.4,-66.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,60.4,-66.2</PageViewport></page 9></circuit>